    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     com.dropbox.attrs    

yJ�rg7�     U(���
